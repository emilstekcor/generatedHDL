-- File Name: reed_solomon/Integer_Output_RS_Decoder_HDL_Optimized.vhd
