module polar_encoder_gamma #(
    parameter int WIDTH = 8
) (
    input  logic signed [WIDTH-1:0] llr_left,
    input  logic signed [WIDTH-1:0] llr_right,
    input  logic u_left,
    output logic signed [WIDTH-1:0] gamma
);
    assign gamma = llr_right + (u_left ? -llr_left : llr_left);
endmodule
